// Code your design here
`include "dat_mem.sv"
`include "top_level_4_260.sv"