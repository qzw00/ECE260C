// Code your testbench here
// or browse Examples
`include "top_tb.sv"